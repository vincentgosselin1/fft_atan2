-- cordic_atan2_v1.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cordic_atan2_v1 is
	port (
		areset : in  std_logic                     := '0';             -- areset.reset
		clk    : in  std_logic                     := '0';             --    clk.clk
		en     : in  std_logic_vector(0 downto 0)  := (others => '0'); --     en.en
		q      : out std_logic_vector(15 downto 0);                    --      q.q
		x      : in  std_logic_vector(15 downto 0) := (others => '0'); --      x.x
		y      : in  std_logic_vector(15 downto 0) := (others => '0')  --      y.y
	);
end entity cordic_atan2_v1;

architecture rtl of cordic_atan2_v1 is
	component cordic_atan2_v1_CORDIC_0 is
		port (
			clk    : in  std_logic                     := 'X';             -- clk
			areset : in  std_logic                     := 'X';             -- reset
			en     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- en
			x      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- x
			y      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- y
			q      : out std_logic_vector(15 downto 0)                     -- q
		);
	end component cordic_atan2_v1_CORDIC_0;

begin

	cordic_0 : component cordic_atan2_v1_CORDIC_0
		port map (
			clk    => clk,    --    clk.clk
			areset => areset, -- areset.reset
			en     => en,     --     en.en
			x      => x,      --      x.x
			y      => y,      --      y.y
			q      => q       --      q.q
		);

end architecture rtl; -- of cordic_atan2_v1
