-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 17.1.0 Build 590 10/25/2017 SJ Lite Edition"
-- CREATED		"Sun Feb 16 12:11:06 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY fft_atan2_v1 IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		RESET :  IN  STD_LOGIC;
		valid :  IN  STD_LOGIC;
		sop :  IN  STD_LOGIC;
		eop :  IN  STD_LOGIC;
		a :  IN  STD_LOGIC;
		b :  IN  STD_LOGIC;
		--real :  IN  STD_LOGIC_VECTOR(15 DOWNTO 0); -- now in the ROM
		c :  OUT  STD_LOGIC;
		rad :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		source_imag :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		source_real :  OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);

		--my additions
		sink_ready : OUT STD_LOGIC;
		mag :  OUT  STD_LOGIC_VECTOR(14 DOWNTO 0);
		source_valid : OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		mag2 : OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		TRIGGER : IN STD_LOGIC--TO START READING ROM.
		
	);
END fft_atan2_v1;

ARCHITECTURE bdf_type OF fft_atan2_v1 IS 

COMPONENT fft_burst_16x1024_v1
	PORT(clk : IN STD_LOGIC;
		 reset_n : IN STD_LOGIC;
		 sink_valid : IN STD_LOGIC;
		 sink_sop : IN STD_LOGIC;
		 sink_eop : IN STD_LOGIC;
		 --inverse : IN STD_LOGIC;
		 inverse : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
		 source_ready : IN STD_LOGIC;
		 sink_error : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 sink_imag : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 sink_real : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 sink_ready : OUT STD_LOGIC;
		 source_valid : OUT STD_LOGIC;
		 source_sop : OUT STD_LOGIC;
		 source_eop : OUT STD_LOGIC;
		 source_error : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		 source_exp : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
		 source_imag : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 source_real : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

--COMPONENT cordic_atan2_v1
--	PORT(areset : IN STD_LOGIC;
--		 clk : IN STD_LOGIC;
--		 en : IN STD_LOGIC;
--		 x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
--		 y : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
--		 q : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
--	);
--END COMPONENT;

--component cordic_atan2_v2 is
--		port (
--			clk    : in  std_logic                     := 'X';             -- clk
--			areset : in  std_logic                     := 'X';             -- reset
--			x      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- x
--			y      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- y
--			q      : out std_logic_vector(15 downto 0);                    -- q
--			r      : out std_logic_vector(15 downto 0);                    -- r
--			en     : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- en
--		);
--	end component cordic_atan2_v2;
	
	component cordic_atan2_v2 is
		port (
			areset : in  std_logic                     := 'X';             -- reset
			clk    : in  std_logic                     := 'X';             -- clk
			en     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- en
			--Angle is q.
			q      : out std_logic_vector(15 downto 0);                    -- q
			--Magnitude is r
			r      : out std_logic_vector(14 downto 0);                    -- r
			x      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- x
			y      : in  std_logic_vector(15 downto 0) := (others => 'X')  -- y
		);
	end component cordic_atan2_v2;
	
component square16bits_v1
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
end component;

component adder32bits_signed
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
end component;

component squareroot32bits_v1
	PORT
	(
		clk		: IN STD_LOGIC ;
		radical		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		q		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		remainder		: OUT STD_LOGIC_VECTOR (16 DOWNTO 0)
	);
end component;

component ROM_RAWDATA
	PORT
	(
		address		: IN STD_LOGIC_VECTOR (9 DOWNTO 0);
		clock		: IN STD_LOGIC  := '1';
		rden		: IN STD_LOGIC  := '1';
		q		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
end component;

COMPONENT ROM_READER_V1
	PORT
	(
		TRIGGER_IN		:	 IN STD_LOGIC;
		CLK		:	 IN STD_LOGIC;
		RESET		:	 IN STD_LOGIC;
		READ_ENA		:	 OUT STD_LOGIC;
		ROM_ADDR		:	 OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;


	

SIGNAL	RESETn :  STD_LOGIC;
SIGNAL	source_imag_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	source_real_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(15 DOWNTO 0);
--SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(0 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(0 TO 1);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(0 DOWNTO 0);
SIGNAL	VCC	:	STD_LOGIC;

SIGNAL	real_sq	: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	imag_sq	: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	w1 : STD_LOGIC;
SIGNAL	dff1 : STD_LOGIC;
SIGNAL	r1	: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL 	remain1	:  STD_LOGIC_VECTOR(16 DOWNTO 0);
SIGNAL	addr : STD_LOGIC_VECTOR (9 DOWNTO 0);
SIGNAL	W3 : STD_LOGIC;
SIGNAL	W4 : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL 	cd1 : STD_LOGIC;
SIGNAL	W5 : STD_LOGIC;
SIGNAL	W6 : STD_LOGIC;




BEGIN 
SYNTHESIZED_WIRE_0 <= "0";
--SYNTHESIZED_WIRE_0 <= '0';
SYNTHESIZED_WIRE_1 <= '1';
SYNTHESIZED_WIRE_2 <= "00";
SYNTHESIZED_WIRE_3 <= "0000000000000000";
VCC <= '1';


--b2v_inst : fft_burst_16x1024_v1
b2v_inst : FFT_Burst_16x1024_v1
PORT MAP(clk => CLK,
		 reset_n => RESETn,
		 sink_valid => valid,
		 sink_sop => sop,
		 sink_eop => eop,
		 inverse => SYNTHESIZED_WIRE_0,
		 source_ready => SYNTHESIZED_WIRE_1,
		 sink_error => SYNTHESIZED_WIRE_2,
		 sink_imag => SYNTHESIZED_WIRE_3,
		 sink_real => W4,
		 source_valid => SYNTHESIZED_WIRE_4(0),
		 source_imag => source_imag_ALTERA_SYNTHESIZED,
		 source_real => source_real_ALTERA_SYNTHESIZED,
		 sink_ready => sink_ready);	


--dff1 data flipflop
process (CLK, RESETn)
begin
	-- Reset whenever the reset signal goes low, regardless of the clock
	-- or the clock enable
	if (RESETn = '0') then
		dff1 <= '0';
	elsif (rising_edge(CLK)) then
			dff1 <= w1;
	end if;
end process;

w1 <= a AND b;
c <= dff1;


--b2v_inst2 : cordic_atan2_v1
--PORT MAP(areset => RESET,
--		 clk => CLK,
--		 en => SYNTHESIZED_WIRE_4(0),
--		 x => source_real_ALTERA_SYNTHESIZED,
--		 y => source_imag_ALTERA_SYNTHESIZED,
--		 q => rad);

	u0 : component cordic_atan2_v2
		port map (
			clk    => CLK,    --    clk.clk
			areset => RESET, -- areset.reset
			x      => source_real_ALTERA_SYNTHESIZED,      --      x.x
			y      => source_imag_ALTERA_SYNTHESIZED,      --      y.y
			q      => rad,      --      q.q
			r      => mag,      --      r.r
			en(0)     => VCC      --     en.en
		);
		
	u1_REAL : component square16bits_v1
		port map (
			clock	=> CLK,
			dataa => source_real_ALTERA_SYNTHESIZED,		
			result => real_sq
		);
		
	u2_IMAG : component square16bits_v1
		port map (
			clock	=> CLK,
			dataa => source_imag_ALTERA_SYNTHESIZED,		
			result => imag_sq
		);
		
	u3: component adder32bits_signed 
	port map
	(
		clock => CLK,
		dataa	=> real_sq,
		datab	=> imag_sq,
		result => r1
	);
	
	u4 : component squareroot32bits_v1
	port map
	(
		clk		=> CLK,
		radical	=> r1,
		q		=> mag2,
		remainder => remain1
	);

	u6 : component ROM_RAWDATA 
	PORT MAP 
	(
		address	 => addr, --output of the counter
		clock	 => CLK,
		rden	 => W6, --activated by count_ena
		q	 => W4
	);
	
	u7 : component ROM_READER_V1
	PORT MAP
	(
		TRIGGER_IN		=> TRIGGER,
		CLK				=> CLK,
		RESET				=> RESET,
		READ_ENA			=> W6,
		ROM_ADDR			=> addr
	);
	
	
	
	
		



		
		

RESETn <= NOT(RESET);
source_valid(0) <= SYNTHESIZED_WIRE_4(0);





source_imag <= source_imag_ALTERA_SYNTHESIZED;
source_real <= source_real_ALTERA_SYNTHESIZED;

END bdf_type;