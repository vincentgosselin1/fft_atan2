// cordic_atan2_v1.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module cordic_atan2_v1 (
		input  wire        areset, // areset.reset
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  en,     //     en.en
		output wire [15:0] q,      //      q.q
		input  wire [15:0] x,      //      x.x
		input  wire [15:0] y       //      y.y
	);

	cordic_atan2_v1_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.en     (en),     //     en.en
		.x      (x),      //      x.x
		.y      (y),      //      y.y
		.q      (q)       //      q.q
	);

endmodule
